module pprows (a, b, c, d, i, o) ;
input a, b, c, d ;
input [15:0] i ;
wire p, q, r, s ;
wire [15:0] w1, w2, w3, w4, w5, w6, w, shift1, shift2, sum, carry ;
output [15:0] o ;

assign p = (~a & ~b & ~c & d) | (~a & ~b & c & ~d) | (a & b & ~c & d) | (a & b & c & ~d) ;
assign q = (~b & c & d) | (b & ~c & ~d) ;
assign r = (~a & b & ~c & d) | (~a & b & c & ~d) | (a & ~b & ~c & d) | (a & ~b & c & ~d) ;
assign s = (~a & b & c & d) | (a & ~b & ~c & ~d) ;

and a1 (w1[15], p, i[15]) ;
and a2 (w1[14], p, i[14]) ;
and a3 (w1[13], p, i[13]) ;
and a4 (w1[12], p, i[12]) ;
and a5 (w1[11], p, i[11]) ;
and a6 (w1[10], p, i[10]) ;
and a7 (w1[9], p, i[9]) ;
and a8 (w1[8], p, i[8]) ;
and a9 (w1[7], p, i[7]) ;
and a10 (w1[6], p, i[6]) ;
and a11 (w1[5], p, i[5]) ;
and a12 (w1[4], p, i[4]) ;
and a13 (w1[3], p, i[3]) ;
and a14 (w1[2], p, i[2]) ;
and a15 (w1[1], p, i[1]) ;
and a16 (w1[0], p, i[0]) ;

buf b1 (shift1[15], i[14]) ;
buf b2 (shift1[14], i[13]) ;
buf b3 (shift1[13], i[12]) ; 
buf b4 (shift1[12], i[11]) ;
buf b5 (shift1[11], i[10]) ;
buf b6 (shift1[10], i[9]) ;
buf b7 (shift1[9], i[8]) ;
buf b8 (shift1[8], i[7]) ;
buf b9 (shift1[7], i[6]) ;
buf b10 (shift1[6], i[5]) ;
buf b11 (shift1[5], i[4]) ;
buf b12 (shift1[4], i[3]) ;
buf b13 (shift1[3], i[2]) ;
buf b14 (shift1[2], i[1]) ;
buf b15 (shift1[1], i[0]) ;
buf b16 (shift1[0], 1'b0) ;

and c1 (w2[15], q, shift1[15]) ;
and c2 (w2[14], q, shift1[14]) ;
and c3 (w2[13], q, shift1[13]) ;
and c4 (w2[12], q, shift1[12]) ;
and c5 (w2[11], q, shift1[11]) ;
and c6 (w2[10], q, shift1[10]) ;
and c7 (w2[9], q, shift1[9]) ;
and c8 (w2[8], q, shift1[8]) ;
and c9 (w2[7], q, shift1[7]) ;
and c10 (w2[6], q, shift1[6]) ;
and c11 (w2[5], q, shift1[5]) ;
and c12 (w2[4], q, shift1[4]) ;
and c13 (w2[3], q, shift1[3]) ;
and c14 (w2[2], q, shift1[2]) ;
and c15 (w2[1], q, shift1[1]) ;
and c16 (w2[0], q, shift1[0]) ;

fa fa1 (i[0], shift1[0], 1'b0, sum[0], carry[0]) ;
fa fa2 (i[1], shift1[1], carry[0], sum[1], carry[1]) ;
fa fa3 (i[2], shift1[2], carry[1], sum[2], carry[2]) ;
fa fa4 (i[3], shift1[3], carry[2], sum[3], carry[3]) ;
fa fa5 (i[4], shift1[4], carry[3], sum[4], carry[4]) ;
fa fa6 (i[5], shift1[5], carry[4], sum[5], carry[5]) ;
fa fa7 (i[6], shift1[6], carry[5], sum[6], carry[6]) ;
fa fa8 (i[7], shift1[7], carry[6], sum[7], carry[7]) ;
fa fa9 (i[8], shift1[8], carry[7], sum[8], carry[8]) ;
fa fa10 (i[9], shift1[9], carry[8], sum[9], carry[9]) ;
fa fa11 (i[10], shift1[10], carry[9], sum[10], carry[10]) ;
fa fa12 (i[11], shift1[11], carry[10], sum[11], carry[11]) ;
fa fa13 (i[12], shift1[12], carry[11], sum[12], carry[12]) ;
fa fa14 (i[13], shift1[13], carry[12], sum[13], carry[13]) ;
fa fa15 (i[14], shift1[14], carry[13], sum[14], carry[14]) ;
fa fa16 (i[15], shift1[15], carry[14], sum[15], carry[15]) ;

and d1 (w3[15], r, sum[15]) ;
and d2 (w3[14], r, sum[14]) ;
and d3 (w3[13], r, sum[13]) ;
and d4 (w3[12], r, sum[12]) ;
and d5 (w3[11], r, sum[11]) ;
and d6 (w3[10], r, sum[10]) ;
and d7 (w3[9], r, sum[9]) ;
and d8 (w3[8], r, sum[8]) ;
and d9 (w3[7], r, sum[7]) ;
and d10 (w3[6], r, sum[6]) ;
and d11 (w3[5], r, sum[5]) ;
and d12 (w3[4], r, sum[4]) ;
and d13 (w3[3], r, sum[3]) ;
and d14 (w3[2], r, sum[2]) ;
and d15 (w3[1], r, sum[1]) ;
and d16 (w3[0], r, sum[0]) ;

buf e1 (shift2[15], shift1[14]) ;
buf e2 (shift2[14], shift1[13]) ;
buf e3 (shift2[13], shift1[12]) ; 
buf e4 (shift2[12], shift1[11]) ;
buf e5 (shift2[11], shift1[10]) ;
buf e6 (shift2[10], shift1[9]) ;
buf e7 (shift2[9], shift1[8]) ;
buf e8 (shift2[8], shift1[7]) ;
buf e9 (shift2[7], shift1[6]) ;
buf e10 (shift2[6], shift1[5]) ;
buf e11 (shift2[5], shift1[4]) ;
buf e12 (shift2[4], shift1[3]) ;
buf e13 (shift2[3], shift1[2]) ;
buf e14 (shift2[2], shift1[1]) ;
buf e15 (shift2[1], shift1[0]) ;
buf e16 (shift2[0], 1'b0) ;

and f1 (w4[15], s, shift2[15]) ;
and f2 (w4[14], s, shift2[14]) ;
and f3 (w4[13], s, shift2[13]) ;
and f4 (w4[12], s, shift2[12]) ;
and f5 (w4[11], s, shift2[11]) ;
and f6 (w4[10], s, shift2[10]) ;
and f7 (w4[9], s, shift2[9]) ;
and f8 (w4[8], s, shift2[8]) ;
and f9 (w4[7], s, shift2[7]) ;
and f10 (w4[6], s, shift2[6]) ;
and f11 (w4[5], s, shift2[5]) ;
and f12 (w4[4], s, shift2[4]) ;
and f13 (w4[3], s, shift2[3]) ;
and f14 (w4[2], s, shift2[2]) ;
and f15 (w4[1], s, shift2[1]) ;
and f16 (w4[0], s, shift2[0]) ;

or g1 (w5[15], w1[15], w2[15]) ;
or g2 (w5[14], w1[14], w2[14]) ;
or g3 (w5[13], w1[13], w2[13]) ;
or g4 (w5[12], w1[12], w2[12]) ;
or g5 (w5[11], w1[11], w2[11]) ;
or g6 (w5[10], w1[10], w2[10]) ;
or g7 (w5[9], w1[9], w2[9]) ;
or g8 (w5[8], w1[8], w2[8]) ;
or g9 (w5[7], w1[7], w2[7]) ;
or g10 (w5[6], w1[6], w2[6]) ;
or g11 (w5[5], w1[5], w2[5]) ;
or g12 (w5[4], w1[4], w2[4]) ;
or g13 (w5[3], w1[3], w2[3]) ;
or g14 (w5[2], w1[2], w2[2]) ;
or g15 (w5[1], w1[1], w2[1]) ;
or g16 (w5[0], w1[0], w2[0]) ;

or h1 (w6[15], w3[15], w4[15]) ;
or h2 (w6[14], w3[14], w4[14]) ;
or h3 (w6[13], w3[13], w4[13]) ;
or h4 (w6[12], w3[12], w4[12]) ;
or h5 (w6[11], w3[11], w4[11]) ;
or h6 (w6[10], w3[10], w4[10]) ;
or h7 (w6[9], w3[9], w4[9]) ;
or h8 (w6[8], w3[8], w4[8]) ;
or h9 (w6[7], w3[7], w4[7]) ;
or h10 (w6[6], w3[6], w4[6]) ;
or h11 (w6[5], w3[5], w4[5]) ;
or h12 (w6[4], w3[4], w4[4]) ;
or h13 (w6[3], w3[3], w4[3]) ;
or h14 (w6[2], w3[2], w4[2]) ;
or h15 (w6[1], w3[1], w4[1]) ;
or h16 (w6[0], w3[0], w4[0]) ;

or j1 (w[15], w5[15], w6[15]) ;
or j2 (w[14], w5[14], w6[14]) ;
or j3 (w[13], w5[13], w6[13]) ;
or j4 (w[12], w5[12], w6[12]) ;
or j5 (w[11], w5[11], w6[11]) ;
or j6 (w[10], w5[10], w6[10]) ;
or j7 (w[9], w5[9], w6[9]) ;
or j8 (w[8], w5[8], w6[8]) ;
or j9 (w[7], w5[7], w6[7]) ;
or j10 (w[6], w5[6], w6[6]) ;
or j11 (w[5], w5[5], w6[5]) ;
or j12 (w[4], w5[4], w6[4]) ;
or j13 (w[3], w5[3], w6[3]) ;
or j14 (w[2], w5[2], w6[2]) ;
or j15 (w[1], w5[1], w6[1]) ;
or j16 (w[0], w5[0], w6[0]) ;

xor k1 (o[15], w[15], a) ;
xor k2 (o[14], w[14], a) ;
xor k3 (o[13], w[13], a) ;
xor k4 (o[12], w[12], a) ;
xor k5 (o[11], w[11], a) ;
xor k6 (o[10], w[10], a) ;
xor k7 (o[9], w[9], a) ;
xor k8 (o[8], w[8], a) ;
xor k9 (o[7], w[7], a) ;
xor k10 (o[6], w[6], a) ;
xor k11 (o[5], w[5], a) ;
xor k12 (o[4], w[4], a) ;
xor k13 (o[3], w[3], a) ;
xor k14 (o[2], w[2], a) ;
xor k15 (o[1], w[1], a) ;
xor k16 (o[0], w[0], a) ;

endmodule
